`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 08/30/2018 10:26:39 AM
// Design Name: 
// Module Name: InstructionMemory_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module InstructionMemory_tb(Instruction);
    reg [31:0] memory;
    output [31:0] Instruction;
    InstructionMemory IM(Address, Instruction);
    
    initial begin
    
        memory[0] = 32'h20100001;	//	main:	addi	$s0, $zero, 1
    memory[1] = 32'h00000000;    //        nop
    memory[2] = 32'h00000000;    //        nop
    memory[3] = 32'h00000000;    //        nop
    memory[4] = 32'h00000000;    //        nop
    memory[5] = 32'h00000000;    //        nop
    memory[6] = 32'h20110001;    //        addi    $s1, $zero, 1
    memory[7] = 32'h00000000;    //        nop
    memory[8] = 32'h00000000;    //        nop
    memory[9] = 32'h00000000;    //        nop
    memory[10] = 32'h00000000;    //        nop
    memory[11] = 32'h00000000;    //        nop
    memory[12] = 32'h02118024;    //        and    $s0, $s0, $s1
    memory[13] = 32'h00000000;    //        nop
    memory[14] = 32'h00000000;    //        nop
    memory[15] = 32'h00000000;    //        nop
    memory[16] = 32'h00000000;    //        nop
    memory[17] = 32'h00000000;    //        nop
    memory[18] = 32'h02008024;    //        and    $s0, $s0, $zero
    memory[19] = 32'h00000000;    //        nop
    memory[20] = 32'h00000000;    //        nop
    memory[21] = 32'h00000000;    //        nop
    memory[22] = 32'h00000000;    //        nop
    memory[23] = 32'h00000000;    //        nop
    memory[24] = 32'h02308022;    //        sub    $s0, $s1, $s0
    memory[25] = 32'h00000000;    //        nop
    memory[26] = 32'h00000000;    //        nop
    memory[27] = 32'h00000000;    //        nop
    memory[28] = 32'h00000000;    //        nop
    memory[29] = 32'h00000000;    //        nop
    memory[30] = 32'h02008027;    //        nor    $s0, $s0, $zero
    memory[31] = 32'h00000000;    //        nop
    memory[32] = 32'h00000000;    //        nop
    memory[33] = 32'h00000000;    //        nop
    memory[34] = 32'h00000000;    //        nop
    memory[35] = 32'h00000000;    //        nop
    memory[36] = 32'h02008027;    //        nor    $s0, $s0, $zero
    memory[37] = 32'h00000000;    //        nop
    memory[38] = 32'h00000000;    //        nop
    memory[39] = 32'h00000000;    //        nop
    memory[40] = 32'h00000000;    //        nop
    memory[41] = 32'h00000000;    //        nop
    memory[42] = 32'h00008025;    //        or    $s0, $zero, $zero
    memory[43] = 32'h00000000;    //        nop
    memory[44] = 32'h00000000;    //        nop
    memory[45] = 32'h00000000;    //        nop
    memory[46] = 32'h00000000;    //        nop
    memory[47] = 32'h00000000;    //        nop
    memory[48] = 32'h02208025;    //        or    $s0, $s1, $zero
    memory[49] = 32'h00000000;    //        nop
    memory[50] = 32'h00000000;    //        nop
    memory[51] = 32'h00000000;    //        nop
    memory[52] = 32'h00000000;    //        nop
    memory[53] = 32'h00000000;    //        nop
    memory[54] = 32'h00108080;    //        sll    $s0, $s0, 2
    memory[55] = 32'h00000000;    //        nop
    memory[56] = 32'h00000000;    //        nop
    memory[57] = 32'h00000000;    //        nop
    memory[58] = 32'h00000000;    //        nop
    memory[59] = 32'h00000000;    //        nop
    memory[60] = 32'h02308004;    //        sllv    $s0, $s0, $s1
    memory[61] = 32'h00000000;    //        nop
    memory[62] = 32'h00000000;    //        nop
    memory[63] = 32'h00000000;    //        nop
    memory[64] = 32'h00000000;    //        nop
    memory[65] = 32'h00000000;    //        nop
    memory[66] = 32'h0200802a;    //        slt    $s0, $s0, $zero
    memory[67] = 32'h00000000;    //        nop
    memory[68] = 32'h00000000;    //        nop
    memory[69] = 32'h00000000;    //        nop
    memory[70] = 32'h00000000;    //        nop
    memory[71] = 32'h00000000;    //        nop
    memory[72] = 32'h0211802a;    //        slt    $s0, $s0, $s1
    memory[73] = 32'h00000000;    //        nop
    memory[74] = 32'h00000000;    //        nop
    memory[75] = 32'h00000000;    //        nop
    memory[76] = 32'h00000000;    //        nop
    memory[77] = 32'h00000000;    //        nop
    memory[78] = 32'h00118043;    //        sra    $s0, $s1, 1
    memory[79] = 32'h00000000;    //        nop
    memory[80] = 32'h00000000;    //        nop
    memory[81] = 32'h00000000;    //        nop
    memory[82] = 32'h00000000;    //        nop
    memory[83] = 32'h00000000;    //        nop
    memory[84] = 32'h00118007;    //        srav    $s0, $s1, $zero
    memory[85] = 32'h00000000;    //        nop
    memory[86] = 32'h00000000;    //        nop
    memory[87] = 32'h00000000;    //        nop
    memory[88] = 32'h00000000;    //        nop
    memory[89] = 32'h00000000;    //        nop
    memory[90] = 32'h00118042;    //        srl    $s0, $s1, 1
    memory[91] = 32'h00000000;    //        nop
    memory[92] = 32'h00000000;    //        nop
    memory[93] = 32'h00000000;    //        nop
    memory[94] = 32'h00000000;    //        nop
    memory[95] = 32'h00000000;    //        nop
    memory[96] = 32'h001180c0;    //        sll    $s0, $s1, 3
    memory[97] = 32'h00000000;    //        nop
    memory[98] = 32'h00000000;    //        nop
    memory[99] = 32'h00000000;    //        nop
    memory[100] = 32'h00000000;    //        nop
    memory[101] = 32'h00000000;    //        nop
    memory[102] = 32'h001080c2;    //        srl    $s0, $s0, 3
    memory[103] = 32'h00000000;    //        nop
    memory[104] = 32'h00000000;    //        nop
    memory[105] = 32'h00000000;    //        nop
    memory[106] = 32'h00000000;    //        nop
    memory[107] = 32'h00000000;    //        nop
    memory[108] = 32'h02308004;    //        sllv    $s0, $s0, $s1
    memory[109] = 32'h00000000;    //        nop
    memory[110] = 32'h00000000;    //        nop
    memory[111] = 32'h00000000;    //        nop
    memory[112] = 32'h00000000;    //        nop
    memory[113] = 32'h00000000;    //        nop
    memory[114] = 32'h02308006;    //        srlv    $s0, $s0, $s1
    memory[115] = 32'h00000000;    //        nop
    memory[116] = 32'h00000000;    //        nop
    memory[117] = 32'h00000000;    //        nop
    memory[118] = 32'h00000000;    //        nop
    memory[119] = 32'h00000000;    //        nop
    memory[120] = 32'h02118026;    //        xor    $s0, $s0, $s1
    memory[121] = 32'h00000000;    //        nop
    memory[122] = 32'h00000000;    //        nop
    memory[123] = 32'h00000000;    //        nop
    memory[124] = 32'h00000000;    //        nop
    memory[125] = 32'h00000000;    //        nop
    memory[126] = 32'h02118026;    //        xor    $s0, $s0, $s1
    memory[127] = 32'h00000000;    //        nop
    memory[128] = 32'h00000000;    //        nop
    memory[129] = 32'h00000000;    //        nop
    memory[130] = 32'h00000000;    //        nop
    memory[131] = 32'h00000000;    //        nop
    memory[132] = 32'h20120004;    //        addi    $s2, $zero, 4
    memory[133] = 32'h00000000;    //        nop
    memory[134] = 32'h00000000;    //        nop
    memory[135] = 32'h00000000;    //        nop
    memory[136] = 32'h00000000;    //        nop
    memory[137] = 32'h00000000;    //        nop
    memory[138] = 32'h72128002;    //        mul    $s0, $s0, $s2
    memory[139] = 32'h00000000;    //        nop
    memory[140] = 32'h00000000;    //        nop
    memory[141] = 32'h00000000;    //        nop
    memory[142] = 32'h00000000;    //        nop
    memory[143] = 32'h00000000;    //        nop
    memory[144] = 32'h22100004;    //        addi    $s0, $s0, 4
    memory[145] = 32'h00000000;    //        nop
    memory[146] = 32'h00000000;    //        nop
    memory[147] = 32'h00000000;    //        nop
    memory[148] = 32'h00000000;    //        nop
    memory[149] = 32'h00000000;    //        nop
    memory[150] = 32'h32100000;    //        andi    $s0, $s0, 0
    memory[151] = 32'h00000000;    //        nop
    memory[152] = 32'h00000000;    //        nop
    memory[153] = 32'h00000000;    //        nop
    memory[154] = 32'h00000000;    //        nop
    memory[155] = 32'h00000000;    //        nop
    memory[156] = 32'h36100001;    //        ori    $s0, $s0, 1
    memory[157] = 32'h00000000;    //        nop
    memory[158] = 32'h00000000;    //        nop
    memory[159] = 32'h00000000;    //        nop
    memory[160] = 32'h00000000;    //        nop
    memory[161] = 32'h00000000;    //        nop
    memory[162] = 32'h2a100000;    //        slti    $s0, $s0, 0
    memory[163] = 32'h00000000;    //        nop
    memory[164] = 32'h00000000;    //        nop
    memory[165] = 32'h00000000;    //        nop
    memory[166] = 32'h00000000;    //        nop
    memory[167] = 32'h00000000;    //        nop
    memory[168] = 32'h2a100001;    //        slti    $s0, $s0, 1
    memory[169] = 32'h00000000;    //        nop
    memory[170] = 32'h00000000;    //        nop
    memory[171] = 32'h00000000;    //        nop
    memory[172] = 32'h00000000;    //        nop
    memory[173] = 32'h00000000;    //        nop
    memory[174] = 32'h3a100001;    //        xori    $s0, $s0, 1
    memory[175] = 32'h00000000;    //        nop
    memory[176] = 32'h00000000;    //        nop
    memory[177] = 32'h00000000;    //        nop
    memory[178] = 32'h00000000;    //        nop
    memory[179] = 32'h00000000;    //        nop
    memory[180] = 32'h3a100001;    //        xori    $s0, $s0, 1
    memory[181] = 32'h00000000;    //        nop
    memory[182] = 32'h00000000;    //        nop
    memory[183] = 32'h00000000;    //        nop
    memory[184] = 32'h00000000;    //        nop
    memory[185] = 32'h00000000;    //        nop
    memory[186] = 32'h2010fffe;    //        addi    $s0, $zero, -2
    memory[187] = 32'h00000000;    //        nop
    memory[188] = 32'h00000000;    //        nop
    memory[189] = 32'h00000000;    //        nop
    memory[190] = 32'h00000000;    //        nop
    memory[191] = 32'h00000000;    //        nop
    memory[192] = 32'h20110002;    //        addi    $s1, $zero, 2
    memory[193] = 32'h00000000;    //        nop
    memory[194] = 32'h00000000;    //        nop
    memory[195] = 32'h00000000;    //        nop
    memory[196] = 32'h00000000;    //        nop
    memory[197] = 32'h00000000;    //        nop
    memory[198] = 32'h0230902b;    //        sltu    $s2, $s1, $s0
    memory[199] = 32'h00000000;    //        nop
    memory[200] = 32'h00000000;    //        nop
    memory[201] = 32'h00000000;    //        nop
    memory[202] = 32'h00000000;    //        nop
    memory[203] = 32'h00000000;    //        nop
    memory[204] = 32'h2e30fffe;    //        sltiu    $s0, $s1, -2
    memory[205] = 32'h00000000;    //        nop
    memory[206] = 32'h00000000;    //        nop
    memory[207] = 32'h00000000;    //        nop
    memory[208] = 32'h00000000;    //        nop
    memory[209] = 32'h00000000;    //        nop
    memory[210] = 32'h0220800a;    //        movz    $s0, $s1, $zero
    memory[211] = 32'h00000000;    //        nop
    memory[212] = 32'h00000000;    //        nop
    memory[213] = 32'h00000000;    //        nop
    memory[214] = 32'h00000000;    //        nop
    memory[215] = 32'h00000000;    //        nop
    memory[216] = 32'h0011800b;    //        movn    $s0, $zero, $s1
    memory[217] = 32'h00000000;    //        nop
    memory[218] = 32'h00000000;    //        nop
    memory[219] = 32'h00000000;    //        nop
    memory[220] = 32'h00000000;    //        nop
    memory[221] = 32'h00000000;    //        nop
    memory[222] = 32'h02328020;    //        add    $s0, $s1, $s2
    memory[223] = 32'h00000000;    //        nop
    memory[224] = 32'h00000000;    //        nop
    memory[225] = 32'h00000000;    //        nop
    memory[226] = 32'h00000000;    //        nop
    memory[227] = 32'h00000000;    //        nop
    memory[228] = 32'h2010fffe;    //        addi    $s0, $zero, -2
    memory[229] = 32'h00000000;    //        nop
    memory[230] = 32'h00000000;    //        nop
    memory[231] = 32'h00000000;    //        nop
    memory[232] = 32'h00000000;    //        nop
    memory[233] = 32'h00000000;    //        nop
    memory[234] = 32'h02308821;    //        addu    $s1, $s1, $s0
    memory[235] = 32'h00000000;    //        nop
    memory[236] = 32'h00000000;    //        nop
    memory[237] = 32'h00000000;    //        nop
    memory[238] = 32'h00000000;    //        nop
    memory[239] = 32'h00000000;    //        nop
    memory[240] = 32'h2411ffff;    //        addiu    $s1, $zero, -1
    memory[241] = 32'h00000000;    //        nop
    memory[242] = 32'h00000000;    //        nop
    memory[243] = 32'h00000000;    //        nop
    memory[244] = 32'h00000000;    //        nop
    memory[245] = 32'h00000000;    //        nop
    memory[246] = 32'h20120020;    //        addi    $s2, $zero, 32
    memory[247] = 32'h00000000;    //        nop
    memory[248] = 32'h00000000;    //        nop
    memory[249] = 32'h00000000;    //        nop
    memory[250] = 32'h00000000;    //        nop
    memory[251] = 32'h00000000;    //        nop
    memory[252] = 32'h02320018;    //        mult    $s1, $s2
    memory[253] = 32'h00000000;    //        nop
    memory[254] = 32'h00000000;    //        nop
    memory[255] = 32'h00000000;    //        nop
    memory[256] = 32'h00000000;    //        nop
    memory[257] = 32'h00000000;    //        nop
    memory[258] = 32'h0000a010;    //        mfhi    $s4
    memory[259] = 32'h00000000;    //        nop
    memory[260] = 32'h00000000;    //        nop
    memory[261] = 32'h00000000;    //        nop
    memory[262] = 32'h00000000;    //        nop
    memory[263] = 32'h00000000;    //        nop
    memory[264] = 32'h0000a812;    //        mflo    $s5
    memory[265] = 32'h00000000;    //        nop
    memory[266] = 32'h00000000;    //        nop
    memory[267] = 32'h00000000;    //        nop
    memory[268] = 32'h00000000;    //        nop
    memory[269] = 32'h00000000;    //        nop
    memory[270] = 32'h02320019;    //        multu    $s1, $s2
    memory[271] = 32'h00000000;    //        nop
    memory[272] = 32'h00000000;    //        nop
    memory[273] = 32'h00000000;    //        nop
    memory[274] = 32'h00000000;    //        nop
    memory[275] = 32'h00000000;    //        nop
    memory[276] = 32'h0000a010;    //        mfhi    $s4
    memory[277] = 32'h00000000;    //        nop
    memory[278] = 32'h00000000;    //        nop
    memory[279] = 32'h00000000;    //        nop
    memory[280] = 32'h00000000;    //        nop
    memory[281] = 32'h00000000;    //        nop
    memory[282] = 32'h0000a812;    //        mflo    $s5
    memory[283] = 32'h00000000;    //        nop
    memory[284] = 32'h00000000;    //        nop
    memory[285] = 32'h00000000;    //        nop
    memory[286] = 32'h00000000;    //        nop
    memory[287] = 32'h00000000;    //        nop
    memory[288] = 32'h72320000;    //        madd    $s1, $s2
    memory[289] = 32'h00000000;    //        nop
    memory[290] = 32'h00000000;    //        nop
    memory[291] = 32'h00000000;    //        nop
    memory[292] = 32'h00000000;    //        nop
    memory[293] = 32'h00000000;    //        nop
    memory[294] = 32'h0000a010;    //        mfhi    $s4
    memory[295] = 32'h00000000;    //        nop
    memory[296] = 32'h00000000;    //        nop
    memory[297] = 32'h00000000;    //        nop
    memory[298] = 32'h00000000;    //        nop
    memory[299] = 32'h00000000;    //        nop
    memory[300] = 32'h0000a812;    //        mflo    $s5
    memory[301] = 32'h00000000;    //        nop
    memory[302] = 32'h00000000;    //        nop
    memory[303] = 32'h00000000;    //        nop
    memory[304] = 32'h00000000;    //        nop
    memory[305] = 32'h00000000;    //        nop
    memory[306] = 32'h02400011;    //        mthi    $s2
    memory[307] = 32'h00000000;    //        nop
    memory[308] = 32'h00000000;    //        nop
    memory[309] = 32'h00000000;    //        nop
    memory[310] = 32'h00000000;    //        nop
    memory[311] = 32'h00000000;    //        nop
    memory[312] = 32'h02200013;    //        mtlo    $s1
    memory[313] = 32'h00000000;    //        nop
    memory[314] = 32'h00000000;    //        nop
    memory[315] = 32'h00000000;    //        nop
    memory[316] = 32'h00000000;    //        nop
    memory[317] = 32'h00000000;    //        nop
    memory[318] = 32'h0000a010;    //        mfhi    $s4
    memory[319] = 32'h00000000;    //        nop
    memory[320] = 32'h00000000;    //        nop
    memory[321] = 32'h00000000;    //        nop
    memory[322] = 32'h00000000;    //        nop
    memory[323] = 32'h00000000;    //        nop
    memory[324] = 32'h0000a812;    //        mflo    $s5
    memory[325] = 32'h00000000;    //        nop
    memory[326] = 32'h00000000;    //        nop
    memory[327] = 32'h00000000;    //        nop
    memory[328] = 32'h00000000;    //        nop
    memory[329] = 32'h00000000;    //        nop
    memory[330] = 32'h3231ffff;    //        andi    $s1, , $s1, 65535
    memory[331] = 32'h00000000;    //        nop
    memory[332] = 32'h00000000;    //        nop
    memory[333] = 32'h00000000;    //        nop
    memory[334] = 32'h00000000;    //        nop
    memory[335] = 32'h00000000;    //        nop
    memory[336] = 32'h72920004;    //        msub    $s4, , $s2
    memory[337] = 32'h00000000;    //        nop
    memory[338] = 32'h00000000;    //        nop
    memory[339] = 32'h00000000;    //        nop
    memory[340] = 32'h00000000;    //        nop
    memory[341] = 32'h00000000;    //        nop
    memory[342] = 32'h0000a010;    //        mfhi    $s4
    memory[343] = 32'h00000000;    //        nop
    memory[344] = 32'h00000000;    //        nop
    memory[345] = 32'h00000000;    //        nop
    memory[346] = 32'h00000000;    //        nop
    memory[347] = 32'h00000000;    //        nop
    memory[348] = 32'h0000a812;    //        mflo    $s5
    memory[349] = 32'h00000000;    //        nop
    memory[350] = 32'h00000000;    //        nop
    memory[351] = 32'h00000000;    //        nop
    memory[352] = 32'h00000000;    //        nop
    memory[353] = 32'h00000000;    //        nop
    memory[354] = 32'h20120001;    //        addi    $s2, $zero, 1
    memory[355] = 32'h00000000;    //        nop
    memory[356] = 32'h00000000;    //        nop
    memory[357] = 32'h00000000;    //        nop
    memory[358] = 32'h00000000;    //        nop
    memory[359] = 32'h00000000;    //        nop
    memory[360] = 32'h00328fc2;    //        rotr    $s1, $s2, 31
    memory[361] = 32'h00000000;    //        nop
    memory[362] = 32'h00000000;    //        nop
    memory[363] = 32'h00000000;    //        nop
    memory[364] = 32'h00000000;    //        nop
    memory[365] = 32'h00000000;    //        nop
    memory[366] = 32'h2014001f;    //        addi    $s4, $zero, 31
    memory[367] = 32'h00000000;    //        nop
    memory[368] = 32'h00000000;    //        nop
    memory[369] = 32'h00000000;    //        nop
    memory[370] = 32'h00000000;    //        nop
    memory[371] = 32'h00000000;    //        nop
    memory[372] = 32'h02918846;    //        rotrv    $s1, $s1, $s4
    memory[373] = 32'h00000000;    //        nop
    memory[374] = 32'h00000000;    //        nop
    memory[375] = 32'h00000000;    //        nop
    memory[376] = 32'h00000000;    //        nop
    memory[377] = 32'h00000000;    //        nop
    memory[378] = 32'h34110ff0;    //        ori    $s1, , $zero, 4080
    memory[379] = 32'h00000000;    //        nop
    memory[380] = 32'h00000000;    //        nop
    memory[381] = 32'h00000000;    //        nop
    memory[382] = 32'h00000000;    //        nop
    memory[383] = 32'h00000000;    //        nop
    memory[384] = 32'h7c11a420;    //        seb    $s4, $s1
    memory[385] = 32'h00000000;    //        nop
    memory[386] = 32'h00000000;    //        nop
    memory[387] = 32'h00000000;    //        nop
    memory[388] = 32'h00000000;    //        nop
    memory[389] = 32'h00000000;    //        nop
    memory[390] = 32'h7c11a620;    //        seh    $s4, , $s1
    memory[391] = 32'h00000000;    //        nop
    memory[392] = 32'h00000000;    //        nop
    memory[393] = 32'h00000000;    //        nop
    memory[394] = 32'h00000000;    //        nop
    memory[395] = 32'h00000000;    //        nop

    end

endmodule
